module adder(input1, input2, out);

       input  [63:0]input1;
       input  [63:0]input2;
       output [63:0]out;


    assign out = input1 + input2; 


endmodule  
